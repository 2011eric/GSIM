module Shreg(out_1, out_2, out_3, out_4, out_5, out_6, in_1, ctrl);
        //parameterize
endmodule